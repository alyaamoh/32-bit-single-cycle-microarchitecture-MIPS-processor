/**************************************************************************************************/
/**************************************************************************************************/
/*****************************		Author: Alyaa Mohamed 	 **************************************/
/*****************************		Module: Shift left twice **************************************/
/**************************************************************************************************/
/**************************************************************************************************/

module shift_left_twice 
#(parameter width=16)
(
    input  wire	[width-1:0] in	,
    
	output reg 	[width-1:0] out
	
);

/***************************************************************************************************/
/***************************************************************************************************/

	always @(*)
		begin
		
			out = in << 2'd2	;
		
		end

endmodule